/*
Copyright (C) 2023, Advanced Micro Devices, Inc. All rights reserved.
SPDX-License-Identifier: MIT
*/


`timescale 1ns / 1ps


module debuglab_top (

);
    
design_1 design_1_i (
);
    
    
endmodule
