// ------------------------------------------------------------------------------
//   (c) Copyright 2020-2021 Advanced Micro Devices, Inc. All rights reserved.
// 
//   This file contains confidential and proprietary information
//   of Advanced Micro Devices, Inc. and is protected under U.S. and
//   international copyright and other intellectual property
//   laws.
// 
//   DISCLAIMER
//   This disclaimer is not a license and does not grant any
//   rights to the materials distributed herewith. Except as
//   otherwise provided in a valid license issued to you by
//   AMD, and to the maximum extent permitted by applicable
//   law: (1) THESE MATERIALS ARE MADE AVAILABLE \"AS IS\" AND
//   WITH ALL FAULTS, AND AMD HEREBY DISCLAIMS ALL WARRANTIES
//   AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
//   BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
//   INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
//   (2) AMD shall not be liable (whether in contract or tort,
//   including negligence, or under any other theory of
//   liability) for any loss or damage of any kind or nature
//   related to, arising under or in connection with these
//   materials, including for any direct, or any indirect,
//   special, incidental, or consequential loss or damage
//   (including loss of data, profits, goodwill, or any type of
//   loss or damage suffered as a result of any action brought
//   by a third party) even if such damage or loss was
//   reasonably foreseeable or AMD had been advised of the
//   possibility of the same.
// 
//   CRITICAL APPLICATIONS
//   AMD products are not designed or intended to be fail-
//   safe, or for use in any application requiring fail-safe
//   performance, such as life-support or safety devices or
//   systems, Class III medical devices, nuclear facilities,
//   applications related to the deployment of airbags, or any
//   other applications that could lead to death, personal
//   injury, or severe property or environmental damage
//   (individually and collectively, \"Critical
//   Applications\"). Customer assumes the sole risk and
//   liability of any use of AMD products in Critical
//   Applications, subject only to applicable laws and
//   regulations governing limitations on product liability.
// 
//   THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
//   PART OF THIS FILE AT ALL TIMES.
// ------------------------------------------------------------------------------
////------------------------------------------------------------------------------


`timescale 1ps/1ps

(* DowngradeIPIdentifiedWarnings="yes" *)
module dcmac_0_prbs_gen_ts (
  clk,
  rst,
  i_id_m1,  // one clock cycle earlier than i_req_num
  i_req_en,
  i_req_num,
  i_seed,
  o_dat
);

  parameter COUNTER_MODE = 0;
  parameter REGISTER_OUTPUT = 1;
  parameter LOAD_SEED = 0;

  input        clk;
  input        rst;
  input        [3-1:0] i_id_m1;
  input        i_req_en;
  input        [8-1:0] i_req_num;
  input        [16-1:0] i_seed;
  output logic [1536-1:0]  o_dat;

  wire   [192+2-1:0][7:0] wide_bus;
  logic  [192:0][2-1:0][7:0] seed_mux;
  logic  [16-1:0] seed_i, seed_o;
  wire   [16-1:0] seed_sel;
  logic  [192-1:0][7:0] cnt_nxt;
  logic  [1536-1:0] prbs_nxt;
  reg    [1536-1:0] dat_reg;
  wire   [1536-1:0] dat_nxt;

  assign dat_nxt = COUNTER_MODE? cnt_nxt : prbs_nxt;
  assign o_dat = REGISTER_OUTPUT? dat_reg : dat_nxt;


  assign wide_bus = {prbs_nxt, seed_o};
  assign seed_i = COUNTER_MODE? {8'd0, cnt_nxt[i_req_num-1]} : seed_mux[i_req_num];
  assign seed_sel = LOAD_SEED? i_seed : seed_o;

  always @* begin
    for (int i=0; i<192; i++) begin
      cnt_nxt[i] = seed_sel + (i + 1);
    end

    for (int i=0; i<=192; i++) begin
      for (int j=0; j<2; j++) begin
        seed_mux[i][j] = wide_bus[i+j];
      end
    end
  end


  always @(posedge clk) begin
    dat_reg <= dat_nxt;
  end

  dcmac_0_ts_context_mem_v2  #(
    .DW (16),
    .INIT_VALUE ({16{1'b1}})
  ) i_dcmac_0_seed_ctx (
    .clk             (clk),
    .rst             (rst),
    .ts_rst          (1'b0),
    .i_rd_id         (i_id_m1),
    .i_ena           (i_req_en),
    .i_dat           (seed_i),
    .o_dat           (seed_o),
    .i_rd_during_wr  (),
    .o_init          ()
  );


  assign prbs_nxt[0] = seed_sel[5]^seed_sel[0]^seed_sel[3]^seed_sel[2];
  assign prbs_nxt[1] = seed_sel[6]^seed_sel[1]^seed_sel[4]^seed_sel[3];
  assign prbs_nxt[2] = seed_sel[4]^seed_sel[5]^seed_sel[7]^seed_sel[2];
  assign prbs_nxt[3] = seed_sel[6]^seed_sel[8]^seed_sel[5]^seed_sel[3];
  assign prbs_nxt[4] = seed_sel[6]^seed_sel[4]^seed_sel[7]^seed_sel[9];
  assign prbs_nxt[5] = seed_sel[10]^seed_sel[8]^seed_sel[5]^seed_sel[7];
  assign prbs_nxt[6] = seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[9];
  assign prbs_nxt[7] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[12];
  assign prbs_nxt[8] = seed_sel[10]^seed_sel[13]^seed_sel[11]^seed_sel[8];
  assign prbs_nxt[9] = seed_sel[14]^seed_sel[11]^seed_sel[9]^seed_sel[12];
  assign prbs_nxt[10] = seed_sel[10]^seed_sel[13]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[11] = seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[5]^seed_sel[3]^seed_sel[0]^seed_sel[2];
  assign prbs_nxt[12] = seed_sel[14]^seed_sel[6]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[3];
  assign prbs_nxt[13] = seed_sel[13]^seed_sel[4]^seed_sel[15]^seed_sel[7]^seed_sel[3]^seed_sel[0];
  assign prbs_nxt[14] = seed_sel[14]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[3]^seed_sel[0]^seed_sel[2];
  assign prbs_nxt[15] = seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[9]^seed_sel[3]^seed_sel[2];
  assign prbs_nxt[16] = seed_sel[6]^seed_sel[10]^seed_sel[4]^seed_sel[0];
  assign prbs_nxt[17] = seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[7];
  assign prbs_nxt[18] = seed_sel[6]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[19] = seed_sel[13]^seed_sel[7]^seed_sel[9]^seed_sel[3];
  assign prbs_nxt[20] = seed_sel[10]^seed_sel[14]^seed_sel[4]^seed_sel[8];
  assign prbs_nxt[21] = seed_sel[11]^seed_sel[5]^seed_sel[9]^seed_sel[15];
  assign prbs_nxt[22] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[23] = seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[4];
  assign prbs_nxt[24] = seed_sel[7]^seed_sel[14]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[25] = seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[26] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[27] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[28] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[29] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[13]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[30] = seed_sel[10]^seed_sel[9]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[31] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[32] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[33] = seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[34] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[35] = seed_sel[10]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[36] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[37] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[38] = seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[1];
  assign prbs_nxt[39] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[14]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[40] = seed_sel[10]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[15];
  assign prbs_nxt[41] = seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[42] = seed_sel[10]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[43] = seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[4];
  assign prbs_nxt[44] = seed_sel[14]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[45] = seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[46] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[47] = seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[48] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[8]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[49] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[13]^seed_sel[8]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[50] = seed_sel[10]^seed_sel[9]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[2];
  assign prbs_nxt[51] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[11]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[52] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[53] = seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[54] = seed_sel[10]^seed_sel[7]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[55] = seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[56] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[57] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[58] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[59] = seed_sel[10]^seed_sel[7]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[60] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[61] = seed_sel[10]^seed_sel[9]^seed_sel[13]^seed_sel[14]^seed_sel[1]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[62] = seed_sel[10]^seed_sel[9]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[63] = seed_sel[10]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[64] = seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[65] = seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[1]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[66] = seed_sel[7]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[8]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[67] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[68] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[69] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[70] = seed_sel[10]^seed_sel[7]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[71] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[72] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[8]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[73] = seed_sel[10]^seed_sel[9]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[74] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[75] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[76] = seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[77] = seed_sel[9]^seed_sel[7]^seed_sel[14]^seed_sel[13]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[78] = seed_sel[10]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[79] = seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[80] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[81] = seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[8];
  assign prbs_nxt[82] = seed_sel[7]^seed_sel[9]^seed_sel[14]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[83] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[84] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[85] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[86] = seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[87] = seed_sel[9]^seed_sel[7]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[88] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[89] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[90] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[91] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[92] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[93] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[94] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[95] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[96] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[97] = seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[98] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[99] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[100] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[101] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[102] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[1];
  assign prbs_nxt[103] = seed_sel[10]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[104] = seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[105] = seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[106] = seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[107] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[108] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[109] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[4];
  assign prbs_nxt[110] = seed_sel[10]^seed_sel[9]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[111] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[112] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[113] = seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[114] = seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[115] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[116] = seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[15];
  assign prbs_nxt[117] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[118] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[119] = seed_sel[7]^seed_sel[9]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[120] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[121] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[122] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[123] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[124] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[125] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[126] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[127] = seed_sel[10]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[128] = seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[129] = seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[130] = seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[131] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[132] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[133] = seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[134] = seed_sel[10]^seed_sel[7]^seed_sel[13]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[135] = seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[136] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[137] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[8]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[138] = seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[2];
  assign prbs_nxt[139] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[140] = seed_sel[10]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[141] = seed_sel[7]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[142] = seed_sel[7]^seed_sel[13]^seed_sel[6]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[143] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[8]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[144] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[1]^seed_sel[8]^seed_sel[15];
  assign prbs_nxt[145] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[146] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[147] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[148] = seed_sel[10]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[149] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[150] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[151] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[152] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[1]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[153] = seed_sel[10]^seed_sel[9]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[154] = seed_sel[10]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[155] = seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[156] = seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[157] = seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[158] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[15];
  assign prbs_nxt[159] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[160] = seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[4];
  assign prbs_nxt[161] = seed_sel[10]^seed_sel[7]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[162] = seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[2];
  assign prbs_nxt[163] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[164] = seed_sel[10]^seed_sel[13]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[165] = seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[2];
  assign prbs_nxt[166] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[167] = seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[8];
  assign prbs_nxt[168] = seed_sel[9]^seed_sel[14]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[169] = seed_sel[10]^seed_sel[13]^seed_sel[6]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[170] = seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[171] = seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[172] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[4]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[173] = seed_sel[10]^seed_sel[9]^seed_sel[14]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[174] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[6]^seed_sel[11]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[175] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[176] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[177] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[14]^seed_sel[13]^seed_sel[4]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[178] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[179] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[180] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[181] = seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[182] = seed_sel[9]^seed_sel[14]^seed_sel[13]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[183] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[184] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[185] = seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[186] = seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[8]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[187] = seed_sel[7]^seed_sel[9]^seed_sel[14]^seed_sel[13]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[2];
  assign prbs_nxt[188] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[189] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[190] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[191] = seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[192] = seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[8]^seed_sel[4]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[193] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[194] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[195] = seed_sel[7]^seed_sel[0]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[196] = seed_sel[0]^seed_sel[13]^seed_sel[1]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[197] = seed_sel[9]^seed_sel[13]^seed_sel[14]^seed_sel[1]^seed_sel[2];
  assign prbs_nxt[198] = seed_sel[10]^seed_sel[3]^seed_sel[14]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[199] = seed_sel[0]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[200] = seed_sel[0]^seed_sel[6]^seed_sel[1]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[201] = seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[1]^seed_sel[2];
  assign prbs_nxt[202] = seed_sel[3]^seed_sel[14]^seed_sel[8]^seed_sel[4]^seed_sel[2];
  assign prbs_nxt[203] = seed_sel[9]^seed_sel[3]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[204] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[4]^seed_sel[2];
  assign prbs_nxt[205] = seed_sel[7]^seed_sel[3]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[206] = seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[207] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[5];
  assign prbs_nxt[208] = seed_sel[10]^seed_sel[7]^seed_sel[14]^seed_sel[6]^seed_sel[4]^seed_sel[8];
  assign prbs_nxt[209] = seed_sel[9]^seed_sel[7]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[210] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[211] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[4];
  assign prbs_nxt[212] = seed_sel[10]^seed_sel[7]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[213] = seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[214] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[215] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[216] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[217] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[218] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[1];
  assign prbs_nxt[219] = seed_sel[10]^seed_sel[9]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[220] = seed_sel[10]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[221] = seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[222] = seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[223] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[8]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[224] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[8]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[225] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[226] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[227] = seed_sel[7]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[228] = seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[229] = seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[230] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[231] = seed_sel[0]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[232] = seed_sel[9]^seed_sel[0]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[233] = seed_sel[10]^seed_sel[13]^seed_sel[1]^seed_sel[2];
  assign prbs_nxt[234] = seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[2];
  assign prbs_nxt[235] = seed_sel[3]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[236] = seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[4]^seed_sel[2];
  assign prbs_nxt[237] = seed_sel[3]^seed_sel[14]^seed_sel[1]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[238] = seed_sel[6]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[239] = seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[2];
  assign prbs_nxt[240] = seed_sel[7]^seed_sel[3]^seed_sel[1]^seed_sel[8];
  assign prbs_nxt[241] = seed_sel[9]^seed_sel[4]^seed_sel[8]^seed_sel[2];
  assign prbs_nxt[242] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[5];
  assign prbs_nxt[243] = seed_sel[10]^seed_sel[6]^seed_sel[11]^seed_sel[4];
  assign prbs_nxt[244] = seed_sel[7]^seed_sel[11]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[245] = seed_sel[13]^seed_sel[6]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[246] = seed_sel[7]^seed_sel[9]^seed_sel[14]^seed_sel[13];
  assign prbs_nxt[247] = seed_sel[10]^seed_sel[14]^seed_sel[8]^seed_sel[15];
  assign prbs_nxt[248] = seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[11]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[249] = seed_sel[10]^seed_sel[0]^seed_sel[6]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[250] = seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[251] = seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[252] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[253] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[2];
  assign prbs_nxt[254] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[255] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[256] = seed_sel[7]^seed_sel[9]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[257] = seed_sel[10]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[258] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[15];
  assign prbs_nxt[259] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[260] = seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[261] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[262] = seed_sel[10]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[263] = seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[264] = seed_sel[10]^seed_sel[6]^seed_sel[13]^seed_sel[1]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[265] = seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[5];
  assign prbs_nxt[266] = seed_sel[6]^seed_sel[14]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[267] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[15];
  assign prbs_nxt[268] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[269] = seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[270] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[271] = seed_sel[7]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[272] = seed_sel[9]^seed_sel[14]^seed_sel[6]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[273] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[15];
  assign prbs_nxt[274] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[275] = seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[276] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[277] = seed_sel[7]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[278] = seed_sel[9]^seed_sel[6]^seed_sel[14]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[279] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[280] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[281] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[282] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[283] = seed_sel[10]^seed_sel[9]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[284] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[285] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[286] = seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[287] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[288] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[289] = seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[290] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[291] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[8];
  assign prbs_nxt[292] = seed_sel[7]^seed_sel[9]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[293] = seed_sel[10]^seed_sel[0]^seed_sel[13]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[294] = seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[295] = seed_sel[10]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[296] = seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[297] = seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[8]^seed_sel[1]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[298] = seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[299] = seed_sel[10]^seed_sel[0]^seed_sel[14]^seed_sel[4];
  assign prbs_nxt[300] = seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[301] = seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[302] = seed_sel[7]^seed_sel[13]^seed_sel[6]^seed_sel[1]^seed_sel[4];
  assign prbs_nxt[303] = seed_sel[7]^seed_sel[14]^seed_sel[8]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[304] = seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[8]^seed_sel[15];
  assign prbs_nxt[305] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[306] = seed_sel[10]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[307] = seed_sel[9]^seed_sel[7]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[308] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[309] = seed_sel[7]^seed_sel[9]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[4];
  assign prbs_nxt[310] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[14]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[311] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[312] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[313] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[314] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[315] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[316] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[317] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[318] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[319] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[320] = seed_sel[10]^seed_sel[9]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[321] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[322] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[323] = seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[324] = seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[1]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[325] = seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[326] = seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[327] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[1]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[328] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[8];
  assign prbs_nxt[329] = seed_sel[9]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[330] = seed_sel[10]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[331] = seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[4];
  assign prbs_nxt[332] = seed_sel[7]^seed_sel[14]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[333] = seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[334] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[335] = seed_sel[10]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[336] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[337] = seed_sel[10]^seed_sel[7]^seed_sel[13]^seed_sel[6]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[338] = seed_sel[7]^seed_sel[9]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[2];
  assign prbs_nxt[339] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[340] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[341] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[342] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[343] = seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[344] = seed_sel[7]^seed_sel[9]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[345] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[346] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[347] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[348] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[1];
  assign prbs_nxt[349] = seed_sel[10]^seed_sel[9]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[350] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[351] = seed_sel[10]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[352] = seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[353] = seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[354] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[355] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[356] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[357] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[358] = seed_sel[10]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[359] = seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[360] = seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[8]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[361] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[8]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[362] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[363] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[11]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[364] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[365] = seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[366] = seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[367] = seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[15];
  assign prbs_nxt[368] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[369] = seed_sel[10]^seed_sel[0]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[370] = seed_sel[9]^seed_sel[0]^seed_sel[11]^seed_sel[1];
  assign prbs_nxt[371] = seed_sel[10]^seed_sel[1]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[372] = seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[2];
  assign prbs_nxt[373] = seed_sel[3]^seed_sel[14]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[374] = seed_sel[13]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[375] = seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[2];
  assign prbs_nxt[376] = seed_sel[7]^seed_sel[3]^seed_sel[4]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[377] = seed_sel[3]^seed_sel[0]^seed_sel[4]^seed_sel[8];
  assign prbs_nxt[378] = seed_sel[9]^seed_sel[4]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[379] = seed_sel[10]^seed_sel[6]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[380] = seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[11];
  assign prbs_nxt[381] = seed_sel[7]^seed_sel[4]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[382] = seed_sel[9]^seed_sel[13]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[383] = seed_sel[10]^seed_sel[9]^seed_sel[6]^seed_sel[14];
  assign prbs_nxt[384] = seed_sel[10]^seed_sel[7]^seed_sel[11]^seed_sel[15];
  assign prbs_nxt[385] = seed_sel[0]^seed_sel[3]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[386] = seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[1]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[387] = seed_sel[10]^seed_sel[7]^seed_sel[14]^seed_sel[13]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[388] = seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[389] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[390] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[2];
  assign prbs_nxt[391] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[392] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[393] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[2];
  assign prbs_nxt[394] = seed_sel[10]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[395] = seed_sel[9]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[396] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[397] = seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[398] = seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[399] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[400] = seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[1];
  assign prbs_nxt[401] = seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[402] = seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[5];
  assign prbs_nxt[403] = seed_sel[10]^seed_sel[7]^seed_sel[14]^seed_sel[6]^seed_sel[1];
  assign prbs_nxt[404] = seed_sel[7]^seed_sel[11]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[405] = seed_sel[9]^seed_sel[0]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[406] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[1];
  assign prbs_nxt[407] = seed_sel[10]^seed_sel[7]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[2];
  assign prbs_nxt[408] = seed_sel[3]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[409] = seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[410] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[1]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[411] = seed_sel[7]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[412] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[413] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[414] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[2];
  assign prbs_nxt[415] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[11]^seed_sel[4]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[416] = seed_sel[10]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[417] = seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[418] = seed_sel[10]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[4]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[419] = seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[420] = seed_sel[0]^seed_sel[14]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[421] = seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[422] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[423] = seed_sel[7]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[424] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[425] = seed_sel[10]^seed_sel[9]^seed_sel[13]^seed_sel[8]^seed_sel[1];
  assign prbs_nxt[426] = seed_sel[10]^seed_sel[9]^seed_sel[14]^seed_sel[11]^seed_sel[2];
  assign prbs_nxt[427] = seed_sel[10]^seed_sel[3]^seed_sel[11]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[428] = seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[429] = seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[430] = seed_sel[7]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[431] = seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[432] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[433] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[1]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[434] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[2];
  assign prbs_nxt[435] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[11]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[436] = seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[437] = seed_sel[10]^seed_sel[9]^seed_sel[13]^seed_sel[14]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[438] = seed_sel[10]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[439] = seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[440] = seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[441] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[1]^seed_sel[8];
  assign prbs_nxt[442] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[14]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[443] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[444] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[445] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[446] = seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[447] = seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[448] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[449] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[450] = seed_sel[9]^seed_sel[0]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[451] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[1]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[452] = seed_sel[10]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[2];
  assign prbs_nxt[453] = seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[454] = seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[455] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[1]^seed_sel[2];
  assign prbs_nxt[456] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[457] = seed_sel[9]^seed_sel[0]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[458] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[1]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[459] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[2];
  assign prbs_nxt[460] = seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[461] = seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[462] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[4]^seed_sel[2];
  assign prbs_nxt[463] = seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[464] = seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[465] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[4]^seed_sel[1]^seed_sel[2];
  assign prbs_nxt[466] = seed_sel[10]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[467] = seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[468] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[4]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[469] = seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[470] = seed_sel[9]^seed_sel[6]^seed_sel[14]^seed_sel[8]^seed_sel[4]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[471] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[472] = seed_sel[10]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[473] = seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[474] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[475] = seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[476] = seed_sel[7]^seed_sel[9]^seed_sel[14]^seed_sel[6]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[477] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[478] = seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[479] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[480] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[481] = seed_sel[9]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[482] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[13]^seed_sel[6]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[483] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[484] = seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[485] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[486] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[2];
  assign prbs_nxt[487] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[488] = seed_sel[10]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[8]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[489] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[2];
  assign prbs_nxt[490] = seed_sel[10]^seed_sel[3]^seed_sel[14]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[491] = seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[492] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[1]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[493] = seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[494] = seed_sel[0]^seed_sel[14]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[495] = seed_sel[13]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[496] = seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[5];
  assign prbs_nxt[497] = seed_sel[7]^seed_sel[6]^seed_sel[1]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[498] = seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[8];
  assign prbs_nxt[499] = seed_sel[9]^seed_sel[8]^seed_sel[4]^seed_sel[1];
  assign prbs_nxt[500] = seed_sel[10]^seed_sel[9]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[501] = seed_sel[10]^seed_sel[3]^seed_sel[6]^seed_sel[11];
  assign prbs_nxt[502] = seed_sel[7]^seed_sel[11]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[503] = seed_sel[13]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[504] = seed_sel[9]^seed_sel[6]^seed_sel[13]^seed_sel[14];
  assign prbs_nxt[505] = seed_sel[10]^seed_sel[7]^seed_sel[14]^seed_sel[15];
  assign prbs_nxt[506] = seed_sel[3]^seed_sel[0]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[507] = seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[508] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[509] = seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[2];
  assign prbs_nxt[510] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[511] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[2];
  assign prbs_nxt[512] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[513] = seed_sel[10]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[514] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[515] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[1]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[516] = seed_sel[9]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[517] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[518] = seed_sel[10]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[519] = seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[520] = seed_sel[7]^seed_sel[13]^seed_sel[6]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[521] = seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[522] = seed_sel[9]^seed_sel[6]^seed_sel[14]^seed_sel[8]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[523] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[524] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[525] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[526] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[527] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[528] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[14]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[529] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[530] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[531] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[532] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[533] = seed_sel[10]^seed_sel[7]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[534] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[535] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[536] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[537] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[538] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[539] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[540] = seed_sel[10]^seed_sel[7]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[541] = seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[542] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[543] = seed_sel[10]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[544] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[545] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[546] = seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[8];
  assign prbs_nxt[547] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[14]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[548] = seed_sel[10]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[549] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[550] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[551] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[552] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[14]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[553] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[15];
  assign prbs_nxt[554] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[555] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[556] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[557] = seed_sel[10]^seed_sel[7]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[558] = seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[559] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[560] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[561] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[562] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[563] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[1];
  assign prbs_nxt[564] = seed_sel[10]^seed_sel[7]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[565] = seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[566] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[567] = seed_sel[10]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[568] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[569] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[8]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[570] = seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[571] = seed_sel[10]^seed_sel[6]^seed_sel[14]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[572] = seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[573] = seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[574] = seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[575] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[576] = seed_sel[10]^seed_sel[7]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[577] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[578] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[13]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[579] = seed_sel[10]^seed_sel[9]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[580] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[581] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[582] = seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[583] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[584] = seed_sel[10]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[585] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[586] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[587] = seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[8];
  assign prbs_nxt[588] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[14]^seed_sel[1]^seed_sel[4]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[589] = seed_sel[10]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[590] = seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[591] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[592] = seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[593] = seed_sel[7]^seed_sel[9]^seed_sel[6]^seed_sel[14]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[594] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[8]^seed_sel[15];
  assign prbs_nxt[595] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[596] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[597] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[598] = seed_sel[10]^seed_sel[7]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[599] = seed_sel[9]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[600] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[601] = seed_sel[10]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[602] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[603] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[604] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[605] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[6]^seed_sel[14]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[606] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[15];
  assign prbs_nxt[607] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[608] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[609] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[610] = seed_sel[10]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[611] = seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[612] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[613] = seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[614] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[615] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[616] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[4];
  assign prbs_nxt[617] = seed_sel[10]^seed_sel[7]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[618] = seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[619] = seed_sel[7]^seed_sel[9]^seed_sel[13]^seed_sel[14]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[620] = seed_sel[10]^seed_sel[13]^seed_sel[14]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[621] = seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[622] = seed_sel[10]^seed_sel[0]^seed_sel[6]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[623] = seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[624] = seed_sel[7]^seed_sel[6]^seed_sel[14]^seed_sel[1]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[625] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[626] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[627] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[628] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[629] = seed_sel[7]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[630] = seed_sel[9]^seed_sel[7]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[631] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[8]^seed_sel[15];
  assign prbs_nxt[632] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[633] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[634] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[635] = seed_sel[10]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[636] = seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[637] = seed_sel[10]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[638] = seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[639] = seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[640] = seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[641] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[1]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[642] = seed_sel[10]^seed_sel[7]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[643] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[8];
  assign prbs_nxt[644] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[8]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[645] = seed_sel[10]^seed_sel[9]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[2];
  assign prbs_nxt[646] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[12];
  assign prbs_nxt[647] = seed_sel[10]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[648] = seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[649] = seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[650] = seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[651] = seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[652] = seed_sel[0]^seed_sel[1]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[653] = seed_sel[0]^seed_sel[3]^seed_sel[1];
  assign prbs_nxt[654] = seed_sel[1]^seed_sel[4]^seed_sel[2];
  assign prbs_nxt[655] = seed_sel[3]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[656] = seed_sel[3]^seed_sel[6]^seed_sel[4];
  assign prbs_nxt[657] = seed_sel[7]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[658] = seed_sel[6]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[659] = seed_sel[7]^seed_sel[9]^seed_sel[6];
  assign prbs_nxt[660] = seed_sel[10]^seed_sel[7]^seed_sel[8];
  assign prbs_nxt[661] = seed_sel[9]^seed_sel[11]^seed_sel[8];
  assign prbs_nxt[662] = seed_sel[10]^seed_sel[9]^seed_sel[12];
  assign prbs_nxt[663] = seed_sel[10]^seed_sel[13]^seed_sel[11];
  assign prbs_nxt[664] = seed_sel[14]^seed_sel[11]^seed_sel[12];
  assign prbs_nxt[665] = seed_sel[13]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[666] = seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[667] = seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[4]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[668] = seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[669] = seed_sel[3]^seed_sel[0]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[2];
  assign prbs_nxt[670] = seed_sel[9]^seed_sel[3]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[671] = seed_sel[10]^seed_sel[3]^seed_sel[6]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[672] = seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[673] = seed_sel[7]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[674] = seed_sel[7]^seed_sel[9]^seed_sel[6]^seed_sel[13]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[675] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[6]^seed_sel[14]^seed_sel[8];
  assign prbs_nxt[676] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[11]^seed_sel[8]^seed_sel[15];
  assign prbs_nxt[677] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[678] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[679] = seed_sel[10]^seed_sel[7]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[680] = seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[681] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[682] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[683] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[15];
  assign prbs_nxt[684] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[685] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[686] = seed_sel[10]^seed_sel[7]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[687] = seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[688] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[689] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[690] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[691] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[692] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[693] = seed_sel[10]^seed_sel[9]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[694] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[695] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[696] = seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[697] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[698] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[699] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[700] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[701] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[8];
  assign prbs_nxt[702] = seed_sel[10]^seed_sel[9]^seed_sel[14]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[703] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[704] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[705] = seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[706] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[707] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[708] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[15];
  assign prbs_nxt[709] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[710] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[711] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[712] = seed_sel[10]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[713] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[714] = seed_sel[10]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[8]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[715] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[716] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[717] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[718] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[719] = seed_sel[9]^seed_sel[7]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[720] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[721] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[722] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[723] = seed_sel[9]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[724] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[12];
  assign prbs_nxt[725] = seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[726] = seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[727] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[728] = seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[4];
  assign prbs_nxt[729] = seed_sel[7]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[730] = seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[731] = seed_sel[7]^seed_sel[9]^seed_sel[14]^seed_sel[6]^seed_sel[1];
  assign prbs_nxt[732] = seed_sel[10]^seed_sel[7]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[733] = seed_sel[9]^seed_sel[0]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[734] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[735] = seed_sel[10]^seed_sel[7]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[2];
  assign prbs_nxt[736] = seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[737] = seed_sel[9]^seed_sel[13]^seed_sel[6]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[738] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[2];
  assign prbs_nxt[739] = seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[15];
  assign prbs_nxt[740] = seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[741] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[1]^seed_sel[4]^seed_sel[2];
  assign prbs_nxt[742] = seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[743] = seed_sel[3]^seed_sel[6]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[744] = seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[4]^seed_sel[2];
  assign prbs_nxt[745] = seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[1]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[746] = seed_sel[9]^seed_sel[6]^seed_sel[8]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[747] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[2];
  assign prbs_nxt[748] = seed_sel[10]^seed_sel[3]^seed_sel[11]^seed_sel[8]^seed_sel[1];
  assign prbs_nxt[749] = seed_sel[9]^seed_sel[11]^seed_sel[4]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[750] = seed_sel[10]^seed_sel[3]^seed_sel[13]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[751] = seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[4];
  assign prbs_nxt[752] = seed_sel[7]^seed_sel[14]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[753] = seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[754] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[755] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[756] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[757] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[6]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[758] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[2];
  assign prbs_nxt[759] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[760] = seed_sel[10]^seed_sel[9]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[761] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[762] = seed_sel[10]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[763] = seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[764] = seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[765] = seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[4]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[766] = seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[767] = seed_sel[0]^seed_sel[3]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[768] = seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[1]^seed_sel[4];
  assign prbs_nxt[769] = seed_sel[7]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[770] = seed_sel[3]^seed_sel[6]^seed_sel[8]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[771] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[4];
  assign prbs_nxt[772] = seed_sel[10]^seed_sel[7]^seed_sel[8]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[773] = seed_sel[9]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[774] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[6]^seed_sel[12];
  assign prbs_nxt[775] = seed_sel[10]^seed_sel[7]^seed_sel[13]^seed_sel[11]^seed_sel[8];
  assign prbs_nxt[776] = seed_sel[9]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[777] = seed_sel[10]^seed_sel[9]^seed_sel[13]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[778] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[779] = seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[780] = seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[781] = seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[2];
  assign prbs_nxt[782] = seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[783] = seed_sel[10]^seed_sel[0]^seed_sel[6]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[784] = seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[11]^seed_sel[1]^seed_sel[2];
  assign prbs_nxt[785] = seed_sel[3]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[786] = seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[787] = seed_sel[10]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[788] = seed_sel[7]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[789] = seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[790] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[8]^seed_sel[1]^seed_sel[4];
  assign prbs_nxt[791] = seed_sel[10]^seed_sel[9]^seed_sel[14]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[792] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[793] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[794] = seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[795] = seed_sel[9]^seed_sel[7]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[796] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[797] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[798] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[799] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[800] = seed_sel[10]^seed_sel[9]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[801] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[802] = seed_sel[10]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[803] = seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[804] = seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[805] = seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[806] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[807] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[808] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[4];
  assign prbs_nxt[809] = seed_sel[10]^seed_sel[9]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[810] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[811] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[812] = seed_sel[7]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[813] = seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[814] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[1]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[815] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[816] = seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[817] = seed_sel[10]^seed_sel[0]^seed_sel[13]^seed_sel[1]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[818] = seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[819] = seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[820] = seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[821] = seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[1]^seed_sel[8]^seed_sel[2];
  assign prbs_nxt[822] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[823] = seed_sel[10]^seed_sel[0]^seed_sel[8]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[824] = seed_sel[9]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[825] = seed_sel[10]^seed_sel[7]^seed_sel[6]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[826] = seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[8];
  assign prbs_nxt[827] = seed_sel[9]^seed_sel[14]^seed_sel[4]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[828] = seed_sel[10]^seed_sel[9]^seed_sel[13]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[829] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[830] = seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[831] = seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[4]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[832] = seed_sel[9]^seed_sel[13]^seed_sel[14]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[833] = seed_sel[10]^seed_sel[9]^seed_sel[14]^seed_sel[6]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[834] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[835] = seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[836] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[1]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[837] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[8]^seed_sel[4]^seed_sel[2];
  assign prbs_nxt[838] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[839] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[840] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[841] = seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[842] = seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[4]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[843] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[844] = seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[845] = seed_sel[9]^seed_sel[0]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[846] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[847] = seed_sel[7]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[2];
  assign prbs_nxt[848] = seed_sel[7]^seed_sel[3]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[849] = seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[850] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[851] = seed_sel[10]^seed_sel[7]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[852] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[11]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[853] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[8]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[854] = seed_sel[10]^seed_sel[9]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[2];
  assign prbs_nxt[855] = seed_sel[10]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[856] = seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[857] = seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[1]^seed_sel[4]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[858] = seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[859] = seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[860] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[861] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[862] = seed_sel[9]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[863] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[864] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4];
  assign prbs_nxt[865] = seed_sel[9]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[866] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[867] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[868] = seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[869] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[870] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[1]^seed_sel[8]^seed_sel[2];
  assign prbs_nxt[871] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[872] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[4]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[873] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[2];
  assign prbs_nxt[874] = seed_sel[10]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[875] = seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[876] = seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[4]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[877] = seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[878] = seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[879] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[880] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[4]^seed_sel[8]^seed_sel[1];
  assign prbs_nxt[881] = seed_sel[9]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[882] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[883] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[4];
  assign prbs_nxt[884] = seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[885] = seed_sel[9]^seed_sel[6]^seed_sel[13]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[886] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[887] = seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[888] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[8]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[889] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[2];
  assign prbs_nxt[890] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[891] = seed_sel[10]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[892] = seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[893] = seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[894] = seed_sel[9]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[4]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[895] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[896] = seed_sel[10]^seed_sel[0]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[897] = seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[898] = seed_sel[10]^seed_sel[7]^seed_sel[6]^seed_sel[13]^seed_sel[1]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[899] = seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[2];
  assign prbs_nxt[900] = seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[4]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[901] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[902] = seed_sel[10]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[2];
  assign prbs_nxt[903] = seed_sel[3]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[904] = seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[905] = seed_sel[7]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[906] = seed_sel[7]^seed_sel[14]^seed_sel[6]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[907] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[908] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[909] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[2];
  assign prbs_nxt[910] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[911] = seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[912] = seed_sel[10]^seed_sel[9]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[913] = seed_sel[10]^seed_sel[7]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[914] = seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[915] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[916] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[8]^seed_sel[1];
  assign prbs_nxt[917] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[918] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[919] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[920] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[921] = seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[922] = seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[8]^seed_sel[4]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[923] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[924] = seed_sel[10]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[925] = seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[926] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[927] = seed_sel[7]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[928] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[929] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[930] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[2];
  assign prbs_nxt[931] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[932] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[933] = seed_sel[10]^seed_sel[9]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[934] = seed_sel[10]^seed_sel[7]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[935] = seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[936] = seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[937] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[938] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[939] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[940] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[941] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[942] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[943] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[944] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[945] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[946] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[947] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[948] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[949] = seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[950] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[951] = seed_sel[10]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[952] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[15];
  assign prbs_nxt[953] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[954] = seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[955] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[6]^seed_sel[14]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[956] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[957] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[958] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[959] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[960] = seed_sel[10]^seed_sel[7]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[961] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[962] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[963] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[964] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[965] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[966] = seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[967] = seed_sel[10]^seed_sel[9]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[968] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[969] = seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[970] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[971] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[1]^seed_sel[8];
  assign prbs_nxt[972] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[973] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[11]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[974] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[975] = seed_sel[10]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[976] = seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[977] = seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[8]^seed_sel[4]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[978] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[979] = seed_sel[10]^seed_sel[0]^seed_sel[14]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[980] = seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[981] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[982] = seed_sel[7]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[983] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[984] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[8]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[985] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[2];
  assign prbs_nxt[986] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[987] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[988] = seed_sel[10]^seed_sel[7]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[989] = seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[990] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[991] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[992] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[993] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[994] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[995] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[996] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[997] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[998] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[999] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1000] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1001] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1002] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1003] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1004] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1005] = seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1006] = seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1007] = seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[1]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[1008] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[1]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[1009] = seed_sel[3]^seed_sel[0]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[1010] = seed_sel[3]^seed_sel[0]^seed_sel[4]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[1011] = seed_sel[13]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1012] = seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1013] = seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[1014] = seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[8]^seed_sel[4]^seed_sel[2];
  assign prbs_nxt[1015] = seed_sel[9]^seed_sel[3]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[1016] = seed_sel[10]^seed_sel[9]^seed_sel[6]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1017] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[5];
  assign prbs_nxt[1018] = seed_sel[7]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[1019] = seed_sel[9]^seed_sel[7]^seed_sel[13]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1020] = seed_sel[10]^seed_sel[9]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[8];
  assign prbs_nxt[1021] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[14]^seed_sel[11]^seed_sel[15];
  assign prbs_nxt[1022] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1023] = seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1024] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1025] = seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1026] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[4]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1027] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1028] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[1029] = seed_sel[10]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1030] = seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1031] = seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[1]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[1032] = seed_sel[9]^seed_sel[7]^seed_sel[13]^seed_sel[14]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1033] = seed_sel[10]^seed_sel[0]^seed_sel[14]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1034] = seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1035] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[1]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1036] = seed_sel[7]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[2];
  assign prbs_nxt[1037] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1038] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[8]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[1039] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[2];
  assign prbs_nxt[1040] = seed_sel[10]^seed_sel[3]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1041] = seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[1042] = seed_sel[7]^seed_sel[14]^seed_sel[13]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1043] = seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1044] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1045] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1046] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[1047] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[6]^seed_sel[8]^seed_sel[1]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1048] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[2];
  assign prbs_nxt[1049] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[1050] = seed_sel[10]^seed_sel[9]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1051] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1052] = seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1053] = seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[8]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1054] = seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1055] = seed_sel[10]^seed_sel[0]^seed_sel[14]^seed_sel[4]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[1056] = seed_sel[3]^seed_sel[0]^seed_sel[11]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[1057] = seed_sel[0]^seed_sel[3]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1058] = seed_sel[13]^seed_sel[6]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1059] = seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1060] = seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[8]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[1061] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[8]^seed_sel[4]^seed_sel[2];
  assign prbs_nxt[1062] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[1063] = seed_sel[10]^seed_sel[9]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1064] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1065] = seed_sel[7]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[1066] = seed_sel[9]^seed_sel[7]^seed_sel[13]^seed_sel[14]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1067] = seed_sel[10]^seed_sel[9]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[8]^seed_sel[15];
  assign prbs_nxt[1068] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1069] = seed_sel[10]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1070] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[1071] = seed_sel[10]^seed_sel[7]^seed_sel[14]^seed_sel[13]^seed_sel[1]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1072] = seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1073] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1074] = seed_sel[10]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1075] = seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1076] = seed_sel[6]^seed_sel[13]^seed_sel[8]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1077] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[5];
  assign prbs_nxt[1078] = seed_sel[10]^seed_sel[6]^seed_sel[14]^seed_sel[8]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[1079] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[11]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1080] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1081] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1082] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1083] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1084] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[8]^seed_sel[4]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1085] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1086] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[1087] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1088] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[1089] = seed_sel[9]^seed_sel[7]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1090] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1091] = seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1092] = seed_sel[10]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1093] = seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[1094] = seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1095] = seed_sel[9]^seed_sel[13]^seed_sel[6]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1096] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[14];
  assign prbs_nxt[1097] = seed_sel[7]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[15];
  assign prbs_nxt[1098] = seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1099] = seed_sel[10]^seed_sel[9]^seed_sel[13]^seed_sel[6]^seed_sel[4]^seed_sel[1];
  assign prbs_nxt[1100] = seed_sel[10]^seed_sel[7]^seed_sel[14]^seed_sel[11]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1101] = seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1102] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1103] = seed_sel[10]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[1104] = seed_sel[9]^seed_sel[7]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1105] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1106] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1107] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[1]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1108] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1109] = seed_sel[10]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1110] = seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1111] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1112] = seed_sel[7]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1113] = seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1114] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1115] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[1]^seed_sel[4]^seed_sel[8];
  assign prbs_nxt[1116] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1117] = seed_sel[10]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1118] = seed_sel[7]^seed_sel[9]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[1119] = seed_sel[10]^seed_sel[7]^seed_sel[14]^seed_sel[13]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1120] = seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[15];
  assign prbs_nxt[1121] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1122] = seed_sel[10]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1123] = seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[1124] = seed_sel[13]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1125] = seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[5];
  assign prbs_nxt[1126] = seed_sel[10]^seed_sel[6]^seed_sel[14]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[1127] = seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[11]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1128] = seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1129] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1130] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1131] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1132] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[8]^seed_sel[4]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1133] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[1134] = seed_sel[10]^seed_sel[9]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1135] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1136] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1137] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1138] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[4]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1139] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1140] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1141] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1142] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1143] = seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1144] = seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1145] = seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1146] = seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1147] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[1148] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[1149] = seed_sel[9]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1150] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1151] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[4];
  assign prbs_nxt[1152] = seed_sel[7]^seed_sel[9]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1153] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1154] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1155] = seed_sel[10]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1156] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1157] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[1]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1158] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1159] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[4]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1160] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1161] = seed_sel[10]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1162] = seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1163] = seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1164] = seed_sel[7]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[1]^seed_sel[8]^seed_sel[15];
  assign prbs_nxt[1165] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1166] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1167] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1];
  assign prbs_nxt[1168] = seed_sel[10]^seed_sel[7]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1169] = seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1170] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[1171] = seed_sel[10]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1172] = seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1173] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1174] = seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[1];
  assign prbs_nxt[1175] = seed_sel[9]^seed_sel[7]^seed_sel[14]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1176] = seed_sel[10]^seed_sel[0]^seed_sel[13]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1177] = seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1178] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1179] = seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4];
  assign prbs_nxt[1180] = seed_sel[9]^seed_sel[14]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1181] = seed_sel[10]^seed_sel[9]^seed_sel[6]^seed_sel[13]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1182] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1183] = seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1184] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1185] = seed_sel[10]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[1186] = seed_sel[7]^seed_sel[9]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1187] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1188] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1189] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[1]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1190] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1191] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1192] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1193] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1194] = seed_sel[7]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1195] = seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1196] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1197] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[1198] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[11]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[1199] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1200] = seed_sel[9]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1201] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1202] = seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[1203] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[8]^seed_sel[4]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1204] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1205] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[1];
  assign prbs_nxt[1206] = seed_sel[10]^seed_sel[11]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1207] = seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1208] = seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[1209] = seed_sel[7]^seed_sel[13]^seed_sel[14]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1210] = seed_sel[0]^seed_sel[14]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1211] = seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1212] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[1213] = seed_sel[7]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[2];
  assign prbs_nxt[1214] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1215] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[4]^seed_sel[8];
  assign prbs_nxt[1216] = seed_sel[10]^seed_sel[9]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[1217] = seed_sel[10]^seed_sel[6]^seed_sel[11]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1218] = seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1219] = seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[1220] = seed_sel[9]^seed_sel[7]^seed_sel[13]^seed_sel[14]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1221] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1222] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1223] = seed_sel[10]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1224] = seed_sel[9]^seed_sel[7]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1225] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1226] = seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[1227] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[4]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1228] = seed_sel[10]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1229] = seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[1230] = seed_sel[13]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1231] = seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[5];
  assign prbs_nxt[1232] = seed_sel[14]^seed_sel[6]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[1233] = seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1234] = seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1235] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1236] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1237] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[1238] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[6]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1239] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[1240] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[1241] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1242] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1243] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1244] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1245] = seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1246] = seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1247] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[1248] = seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1249] = seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1250] = seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[1]^seed_sel[4];
  assign prbs_nxt[1251] = seed_sel[14]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1252] = seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1253] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1254] = seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[1255] = seed_sel[9]^seed_sel[7]^seed_sel[6]^seed_sel[8]^seed_sel[4]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1256] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[1257] = seed_sel[10]^seed_sel[9]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[4];
  assign prbs_nxt[1258] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[11]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1259] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1260] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[1261] = seed_sel[10]^seed_sel[7]^seed_sel[13]^seed_sel[14]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1262] = seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1263] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1264] = seed_sel[10]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1265] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1266] = seed_sel[10]^seed_sel[7]^seed_sel[13]^seed_sel[6]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1267] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8];
  assign prbs_nxt[1268] = seed_sel[10]^seed_sel[9]^seed_sel[14]^seed_sel[1]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1269] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1270] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1271] = seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1272] = seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[8]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[1273] = seed_sel[9]^seed_sel[7]^seed_sel[14]^seed_sel[13]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1274] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1275] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1276] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[1277] = seed_sel[7]^seed_sel[9]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1278] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1279] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[1280] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1281] = seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1282] = seed_sel[10]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[1283] = seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1284] = seed_sel[0]^seed_sel[14]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1285] = seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1286] = seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[4]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[1287] = seed_sel[7]^seed_sel[6]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1288] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[1289] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[6]^seed_sel[1]^seed_sel[8];
  assign prbs_nxt[1290] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[11]^seed_sel[8]^seed_sel[2];
  assign prbs_nxt[1291] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[11]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[1292] = seed_sel[10]^seed_sel[9]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[1293] = seed_sel[10]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1294] = seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1295] = seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1296] = seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1297] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[1298] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1299] = seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[1300] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[6]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1301] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1302] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[1303] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[13]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1304] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[2];
  assign prbs_nxt[1305] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1306] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1307] = seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1308] = seed_sel[10]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[4]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1309] = seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[1310] = seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1311] = seed_sel[0]^seed_sel[13]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1312] = seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[1];
  assign prbs_nxt[1313] = seed_sel[10]^seed_sel[7]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1314] = seed_sel[0]^seed_sel[11]^seed_sel[8];
  assign prbs_nxt[1315] = seed_sel[9]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[1316] = seed_sel[10]^seed_sel[13]^seed_sel[2];
  assign prbs_nxt[1317] = seed_sel[3]^seed_sel[14]^seed_sel[11];
  assign prbs_nxt[1318] = seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1319] = seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[2];
  assign prbs_nxt[1320] = seed_sel[3]^seed_sel[14]^seed_sel[4]^seed_sel[1];
  assign prbs_nxt[1321] = seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1322] = seed_sel[0]^seed_sel[6]^seed_sel[2];
  assign prbs_nxt[1323] = seed_sel[7]^seed_sel[3]^seed_sel[1];
  assign prbs_nxt[1324] = seed_sel[4]^seed_sel[8]^seed_sel[2];
  assign prbs_nxt[1325] = seed_sel[9]^seed_sel[3]^seed_sel[5];
  assign prbs_nxt[1326] = seed_sel[10]^seed_sel[6]^seed_sel[4];
  assign prbs_nxt[1327] = seed_sel[7]^seed_sel[11]^seed_sel[5];
  assign prbs_nxt[1328] = seed_sel[6]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[1329] = seed_sel[7]^seed_sel[9]^seed_sel[13];
  assign prbs_nxt[1330] = seed_sel[10]^seed_sel[14]^seed_sel[8];
  assign prbs_nxt[1331] = seed_sel[9]^seed_sel[11]^seed_sel[15];
  assign prbs_nxt[1332] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1333] = seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[4];
  assign prbs_nxt[1334] = seed_sel[7]^seed_sel[14]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1335] = seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1336] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1337] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1338] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[4];
  assign prbs_nxt[1339] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1340] = seed_sel[10]^seed_sel[9]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1341] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[12];
  assign prbs_nxt[1342] = seed_sel[10]^seed_sel[7]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1343] = seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1344] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1345] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[1346] = seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1347] = seed_sel[0]^seed_sel[13]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1348] = seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[1];
  assign prbs_nxt[1349] = seed_sel[14]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1350] = seed_sel[0]^seed_sel[15];
  assign prbs_nxt[1351] = seed_sel[3]^seed_sel[0]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1352] = seed_sel[3]^seed_sel[6]^seed_sel[4]^seed_sel[1]^seed_sel[2];
  assign prbs_nxt[1353] = seed_sel[7]^seed_sel[3]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1354] = seed_sel[3]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[1355] = seed_sel[9]^seed_sel[7]^seed_sel[6]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[1356] = seed_sel[10]^seed_sel[7]^seed_sel[6]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[1357] = seed_sel[7]^seed_sel[9]^seed_sel[6]^seed_sel[11]^seed_sel[8];
  assign prbs_nxt[1358] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[1359] = seed_sel[10]^seed_sel[9]^seed_sel[13]^seed_sel[11]^seed_sel[8];
  assign prbs_nxt[1360] = seed_sel[10]^seed_sel[9]^seed_sel[14]^seed_sel[11]^seed_sel[12];
  assign prbs_nxt[1361] = seed_sel[10]^seed_sel[13]^seed_sel[11]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1362] = seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1363] = seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1364] = seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[1365] = seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1366] = seed_sel[9]^seed_sel[0]^seed_sel[1]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[1367] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[1];
  assign prbs_nxt[1368] = seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[2];
  assign prbs_nxt[1369] = seed_sel[3]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1370] = seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[4];
  assign prbs_nxt[1371] = seed_sel[7]^seed_sel[14]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[1372] = seed_sel[6]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1373] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1374] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[8]^seed_sel[4]^seed_sel[1];
  assign prbs_nxt[1375] = seed_sel[9]^seed_sel[7]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1376] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1377] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[4];
  assign prbs_nxt[1378] = seed_sel[10]^seed_sel[7]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1379] = seed_sel[9]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1380] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1381] = seed_sel[10]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[1382] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1383] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1384] = seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[1];
  assign prbs_nxt[1385] = seed_sel[10]^seed_sel[14]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1386] = seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1387] = seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1388] = seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1389] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[4]^seed_sel[8];
  assign prbs_nxt[1390] = seed_sel[10]^seed_sel[9]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1391] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[5];
  assign prbs_nxt[1392] = seed_sel[10]^seed_sel[7]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[1393] = seed_sel[7]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1394] = seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[1395] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[13]^seed_sel[14]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[1396] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1397] = seed_sel[9]^seed_sel[0]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1398] = seed_sel[10]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[1399] = seed_sel[7]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[2];
  assign prbs_nxt[1400] = seed_sel[3]^seed_sel[14]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1401] = seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1402] = seed_sel[10]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[1]^seed_sel[2];
  assign prbs_nxt[1403] = seed_sel[7]^seed_sel[3]^seed_sel[11]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1404] = seed_sel[0]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1405] = seed_sel[9]^seed_sel[6]^seed_sel[13]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[1406] = seed_sel[10]^seed_sel[7]^seed_sel[6]^seed_sel[14]^seed_sel[2];
  assign prbs_nxt[1407] = seed_sel[7]^seed_sel[3]^seed_sel[11]^seed_sel[8]^seed_sel[15];
  assign prbs_nxt[1408] = seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1409] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[4]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[1410] = seed_sel[10]^seed_sel[7]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1411] = seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1412] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1413] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[1414] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1415] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1416] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1417] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1418] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1419] = seed_sel[10]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1420] = seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1421] = seed_sel[10]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1422] = seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1423] = seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1424] = seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[1425] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[1]^seed_sel[4]^seed_sel[8];
  assign prbs_nxt[1426] = seed_sel[10]^seed_sel[9]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1427] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[11];
  assign prbs_nxt[1428] = seed_sel[10]^seed_sel[7]^seed_sel[11]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[1429] = seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1430] = seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[12];
  assign prbs_nxt[1431] = seed_sel[10]^seed_sel[14]^seed_sel[13]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[1432] = seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1433] = seed_sel[0]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1434] = seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[1];
  assign prbs_nxt[1435] = seed_sel[7]^seed_sel[14]^seed_sel[1]^seed_sel[2];
  assign prbs_nxt[1436] = seed_sel[3]^seed_sel[8]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1437] = seed_sel[9]^seed_sel[0]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1438] = seed_sel[10]^seed_sel[3]^seed_sel[6]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[1439] = seed_sel[7]^seed_sel[6]^seed_sel[11]^seed_sel[4]^seed_sel[2];
  assign prbs_nxt[1440] = seed_sel[7]^seed_sel[3]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1441] = seed_sel[9]^seed_sel[6]^seed_sel[13]^seed_sel[8]^seed_sel[4];
  assign prbs_nxt[1442] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[14]^seed_sel[5];
  assign prbs_nxt[1443] = seed_sel[10]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[15];
  assign prbs_nxt[1444] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[11]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1445] = seed_sel[10]^seed_sel[3]^seed_sel[13]^seed_sel[6]^seed_sel[8]^seed_sel[4]^seed_sel[1]^seed_sel[12];
  assign prbs_nxt[1446] = seed_sel[9]^seed_sel[7]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1447] = seed_sel[10]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1448] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1449] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[4]^seed_sel[1]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1450] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1451] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1452] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1453] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1454] = seed_sel[7]^seed_sel[9]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1455] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[1456] = seed_sel[10]^seed_sel[9]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[1457] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1458] = seed_sel[10]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1459] = seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[1460] = seed_sel[7]^seed_sel[14]^seed_sel[13]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1461] = seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1462] = seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1463] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[6]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1464] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[1];
  assign prbs_nxt[1465] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[8]^seed_sel[1]^seed_sel[4]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1466] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1467] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[1468] = seed_sel[10]^seed_sel[7]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1469] = seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1470] = seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1471] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[8]^seed_sel[4]^seed_sel[15];
  assign prbs_nxt[1472] = seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1473] = seed_sel[10]^seed_sel[0]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1474] = seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[1];
  assign prbs_nxt[1475] = seed_sel[14]^seed_sel[4]^seed_sel[1]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1476] = seed_sel[3]^seed_sel[13]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1477] = seed_sel[0]^seed_sel[14]^seed_sel[6]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1478] = seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1479] = seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[5];
  assign prbs_nxt[1480] = seed_sel[7]^seed_sel[9]^seed_sel[6]^seed_sel[1]^seed_sel[8]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[1481] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[6]^seed_sel[8]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1482] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[8];
  assign prbs_nxt[1483] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[12];
  assign prbs_nxt[1484] = seed_sel[10]^seed_sel[9]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1485] = seed_sel[10]^seed_sel[9]^seed_sel[13]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[12];
  assign prbs_nxt[1486] = seed_sel[10]^seed_sel[7]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1487] = seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1488] = seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1489] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[1]^seed_sel[15];
  assign prbs_nxt[1490] = seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1491] = seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1492] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[6]^seed_sel[1]^seed_sel[4];
  assign prbs_nxt[1493] = seed_sel[10]^seed_sel[7]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1494] = seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1495] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[4]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1496] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5];
  assign prbs_nxt[1497] = seed_sel[7]^seed_sel[9]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1498] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[0]^seed_sel[13]^seed_sel[8]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1499] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1500] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1501] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[13]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1502] = seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[1]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1503] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[1]^seed_sel[4]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1504] = seed_sel[10]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[4]^seed_sel[8]^seed_sel[15];
  assign prbs_nxt[1505] = seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[11]^seed_sel[1]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1506] = seed_sel[10]^seed_sel[0]^seed_sel[1]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1507] = seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[1];
  assign prbs_nxt[1508] = seed_sel[7]^seed_sel[14]^seed_sel[4]^seed_sel[1]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1509] = seed_sel[3]^seed_sel[13]^seed_sel[8]^seed_sel[5]^seed_sel[15]^seed_sel[2];
  assign prbs_nxt[1510] = seed_sel[9]^seed_sel[0]^seed_sel[6]^seed_sel[14]^seed_sel[4]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1511] = seed_sel[10]^seed_sel[7]^seed_sel[3]^seed_sel[6]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1512] = seed_sel[7]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5];
  assign prbs_nxt[1513] = seed_sel[9]^seed_sel[7]^seed_sel[6]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[12];
  assign prbs_nxt[1514] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[13]^seed_sel[6]^seed_sel[8]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1515] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[3]^seed_sel[14]^seed_sel[6]^seed_sel[11]^seed_sel[8];
  assign prbs_nxt[1516] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1517] = seed_sel[10]^seed_sel[9]^seed_sel[0]^seed_sel[3]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1518] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[1]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[1519] = seed_sel[10]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1520] = seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[11]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1521] = seed_sel[7]^seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[1]^seed_sel[5]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1522] = seed_sel[0]^seed_sel[14]^seed_sel[13]^seed_sel[6]^seed_sel[1]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1523] = seed_sel[9]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[1]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1524] = seed_sel[10]^seed_sel[7]^seed_sel[0]^seed_sel[3]^seed_sel[6]^seed_sel[1]^seed_sel[4]^seed_sel[8]^seed_sel[5]^seed_sel[15];
  assign prbs_nxt[1525] = seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[11]^seed_sel[8]^seed_sel[1]^seed_sel[4];
  assign prbs_nxt[1526] = seed_sel[10]^seed_sel[9]^seed_sel[7]^seed_sel[4]^seed_sel[8]^seed_sel[1]^seed_sel[5]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1527] = seed_sel[10]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[5]^seed_sel[2];
  assign prbs_nxt[1528] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[6]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[12];
  assign prbs_nxt[1529] = seed_sel[10]^seed_sel[7]^seed_sel[13]^seed_sel[11]^seed_sel[8]^seed_sel[4]^seed_sel[5]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1530] = seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[6]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[8]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1531] = seed_sel[10]^seed_sel[7]^seed_sel[9]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1532] = seed_sel[10]^seed_sel[3]^seed_sel[0]^seed_sel[13]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[8]^seed_sel[15];
  assign prbs_nxt[1533] = seed_sel[9]^seed_sel[3]^seed_sel[0]^seed_sel[14]^seed_sel[11]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12]^seed_sel[2];
  assign prbs_nxt[1534] = seed_sel[10]^seed_sel[0]^seed_sel[13]^seed_sel[4]^seed_sel[1]^seed_sel[15]^seed_sel[12];
  assign prbs_nxt[1535] = seed_sel[0]^seed_sel[3]^seed_sel[14]^seed_sel[13]^seed_sel[11]^seed_sel[1];

endmodule
